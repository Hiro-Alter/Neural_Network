// RedNeuronal_NiosII_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module RedNeuronal_NiosII_tb (
	);

	wire    redneuronal_niosii_inst_clk_bfm_clk_clk; // RedNeuronal_NiosII_inst_clk_bfm:clk -> RedNeuronal_NiosII_inst:clk_clk

	RedNeuronal_NiosII redneuronal_niosii_inst (
		.clk_clk (redneuronal_niosii_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) redneuronal_niosii_inst_clk_bfm (
		.clk (redneuronal_niosii_inst_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
