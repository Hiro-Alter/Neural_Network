// RedNeuronal_NiosII.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module RedNeuronal_NiosII (
		input  wire  clk_clk  // clk.clk
	);

	wire         redneuronal_niosii_debug_reset_request_reset;                     // RedNeuronal_NiosII:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] redneuronal_niosii_data_master_readdata;                          // mm_interconnect_0:RedNeuronal_NiosII_data_master_readdata -> RedNeuronal_NiosII:d_readdata
	wire         redneuronal_niosii_data_master_waitrequest;                       // mm_interconnect_0:RedNeuronal_NiosII_data_master_waitrequest -> RedNeuronal_NiosII:d_waitrequest
	wire         redneuronal_niosii_data_master_debugaccess;                       // RedNeuronal_NiosII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:RedNeuronal_NiosII_data_master_debugaccess
	wire  [20:0] redneuronal_niosii_data_master_address;                           // RedNeuronal_NiosII:d_address -> mm_interconnect_0:RedNeuronal_NiosII_data_master_address
	wire   [3:0] redneuronal_niosii_data_master_byteenable;                        // RedNeuronal_NiosII:d_byteenable -> mm_interconnect_0:RedNeuronal_NiosII_data_master_byteenable
	wire         redneuronal_niosii_data_master_read;                              // RedNeuronal_NiosII:d_read -> mm_interconnect_0:RedNeuronal_NiosII_data_master_read
	wire         redneuronal_niosii_data_master_write;                             // RedNeuronal_NiosII:d_write -> mm_interconnect_0:RedNeuronal_NiosII_data_master_write
	wire  [31:0] redneuronal_niosii_data_master_writedata;                         // RedNeuronal_NiosII:d_writedata -> mm_interconnect_0:RedNeuronal_NiosII_data_master_writedata
	wire  [31:0] redneuronal_niosii_instruction_master_readdata;                   // mm_interconnect_0:RedNeuronal_NiosII_instruction_master_readdata -> RedNeuronal_NiosII:i_readdata
	wire         redneuronal_niosii_instruction_master_waitrequest;                // mm_interconnect_0:RedNeuronal_NiosII_instruction_master_waitrequest -> RedNeuronal_NiosII:i_waitrequest
	wire  [20:0] redneuronal_niosii_instruction_master_address;                    // RedNeuronal_NiosII:i_address -> mm_interconnect_0:RedNeuronal_NiosII_instruction_master_address
	wire         redneuronal_niosii_instruction_master_read;                       // RedNeuronal_NiosII:i_read -> mm_interconnect_0:RedNeuronal_NiosII_instruction_master_read
	wire         mm_interconnect_0_uart_avalon_jtag_slave_chipselect;              // mm_interconnect_0:uart_avalon_jtag_slave_chipselect -> uart:av_chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_readdata;                // uart:av_readdata -> mm_interconnect_0:uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_waitrequest;             // uart:av_waitrequest -> mm_interconnect_0:uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart_avalon_jtag_slave_address;                 // mm_interconnect_0:uart_avalon_jtag_slave_address -> uart:av_address
	wire         mm_interconnect_0_uart_avalon_jtag_slave_read;                    // mm_interconnect_0:uart_avalon_jtag_slave_read -> uart:av_read_n
	wire         mm_interconnect_0_uart_avalon_jtag_slave_write;                   // mm_interconnect_0:uart_avalon_jtag_slave_write -> uart:av_write_n
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_writedata;               // mm_interconnect_0:uart_avalon_jtag_slave_writedata -> uart:av_writedata
	wire  [31:0] mm_interconnect_0_redneuronal_niosii_debug_mem_slave_readdata;    // RedNeuronal_NiosII:debug_mem_slave_readdata -> mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_readdata
	wire         mm_interconnect_0_redneuronal_niosii_debug_mem_slave_waitrequest; // RedNeuronal_NiosII:debug_mem_slave_waitrequest -> mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_redneuronal_niosii_debug_mem_slave_debugaccess; // mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_debugaccess -> RedNeuronal_NiosII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_redneuronal_niosii_debug_mem_slave_address;     // mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_address -> RedNeuronal_NiosII:debug_mem_slave_address
	wire         mm_interconnect_0_redneuronal_niosii_debug_mem_slave_read;        // mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_read -> RedNeuronal_NiosII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_redneuronal_niosii_debug_mem_slave_byteenable;  // mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_byteenable -> RedNeuronal_NiosII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_redneuronal_niosii_debug_mem_slave_write;       // mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_write -> RedNeuronal_NiosII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_redneuronal_niosii_debug_mem_slave_writedata;   // mm_interconnect_0:RedNeuronal_NiosII_debug_mem_slave_writedata -> RedNeuronal_NiosII:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                             // mm_interconnect_0:sram_s1_chipselect -> sram:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                               // sram:readdata -> mm_interconnect_0:sram_s1_readdata
	wire  [16:0] mm_interconnect_0_sram_s1_address;                                // mm_interconnect_0:sram_s1_address -> sram:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                             // mm_interconnect_0:sram_s1_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_s1_write;                                  // mm_interconnect_0:sram_s1_write -> sram:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                              // mm_interconnect_0:sram_s1_writedata -> sram:writedata
	wire         mm_interconnect_0_sram_s1_clken;                                  // mm_interconnect_0:sram_s1_clken -> sram:clken
	wire         irq_mapper_receiver0_irq;                                         // uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] redneuronal_niosii_irq_irq;                                       // irq_mapper:sender_irq -> RedNeuronal_NiosII:irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [RedNeuronal_NiosII:reset_n, irq_mapper:reset, mm_interconnect_0:RedNeuronal_NiosII_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sram:reset, uart:rst_n]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [RedNeuronal_NiosII:reset_req, rst_translator:reset_req_in, sram:reset_req]

	RedNeuronal_NiosII_RedNeuronal_NiosII redneuronal_niosii (
		.clk                                 (clk_clk),                                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                                  //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                               //                          .reset_req
		.d_address                           (redneuronal_niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (redneuronal_niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (redneuronal_niosii_data_master_read),                              //                          .read
		.d_readdata                          (redneuronal_niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (redneuronal_niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (redneuronal_niosii_data_master_write),                             //                          .write
		.d_writedata                         (redneuronal_niosii_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (redneuronal_niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (redneuronal_niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (redneuronal_niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (redneuronal_niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (redneuronal_niosii_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (redneuronal_niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (redneuronal_niosii_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                                  // custom_instruction_master.readra
	);

	RedNeuronal_NiosII_sram sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	RedNeuronal_NiosII_uart uart (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	RedNeuronal_NiosII_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                        (clk_clk),                                                          //                                      clk_0_clk.clk
		.RedNeuronal_NiosII_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                   // RedNeuronal_NiosII_reset_reset_bridge_in_reset.reset
		.RedNeuronal_NiosII_data_master_address               (redneuronal_niosii_data_master_address),                           //                 RedNeuronal_NiosII_data_master.address
		.RedNeuronal_NiosII_data_master_waitrequest           (redneuronal_niosii_data_master_waitrequest),                       //                                               .waitrequest
		.RedNeuronal_NiosII_data_master_byteenable            (redneuronal_niosii_data_master_byteenable),                        //                                               .byteenable
		.RedNeuronal_NiosII_data_master_read                  (redneuronal_niosii_data_master_read),                              //                                               .read
		.RedNeuronal_NiosII_data_master_readdata              (redneuronal_niosii_data_master_readdata),                          //                                               .readdata
		.RedNeuronal_NiosII_data_master_write                 (redneuronal_niosii_data_master_write),                             //                                               .write
		.RedNeuronal_NiosII_data_master_writedata             (redneuronal_niosii_data_master_writedata),                         //                                               .writedata
		.RedNeuronal_NiosII_data_master_debugaccess           (redneuronal_niosii_data_master_debugaccess),                       //                                               .debugaccess
		.RedNeuronal_NiosII_instruction_master_address        (redneuronal_niosii_instruction_master_address),                    //          RedNeuronal_NiosII_instruction_master.address
		.RedNeuronal_NiosII_instruction_master_waitrequest    (redneuronal_niosii_instruction_master_waitrequest),                //                                               .waitrequest
		.RedNeuronal_NiosII_instruction_master_read           (redneuronal_niosii_instruction_master_read),                       //                                               .read
		.RedNeuronal_NiosII_instruction_master_readdata       (redneuronal_niosii_instruction_master_readdata),                   //                                               .readdata
		.RedNeuronal_NiosII_debug_mem_slave_address           (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_address),     //             RedNeuronal_NiosII_debug_mem_slave.address
		.RedNeuronal_NiosII_debug_mem_slave_write             (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_write),       //                                               .write
		.RedNeuronal_NiosII_debug_mem_slave_read              (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_read),        //                                               .read
		.RedNeuronal_NiosII_debug_mem_slave_readdata          (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_readdata),    //                                               .readdata
		.RedNeuronal_NiosII_debug_mem_slave_writedata         (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_writedata),   //                                               .writedata
		.RedNeuronal_NiosII_debug_mem_slave_byteenable        (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_byteenable),  //                                               .byteenable
		.RedNeuronal_NiosII_debug_mem_slave_waitrequest       (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_waitrequest), //                                               .waitrequest
		.RedNeuronal_NiosII_debug_mem_slave_debugaccess       (mm_interconnect_0_redneuronal_niosii_debug_mem_slave_debugaccess), //                                               .debugaccess
		.sram_s1_address                                      (mm_interconnect_0_sram_s1_address),                                //                                        sram_s1.address
		.sram_s1_write                                        (mm_interconnect_0_sram_s1_write),                                  //                                               .write
		.sram_s1_readdata                                     (mm_interconnect_0_sram_s1_readdata),                               //                                               .readdata
		.sram_s1_writedata                                    (mm_interconnect_0_sram_s1_writedata),                              //                                               .writedata
		.sram_s1_byteenable                                   (mm_interconnect_0_sram_s1_byteenable),                             //                                               .byteenable
		.sram_s1_chipselect                                   (mm_interconnect_0_sram_s1_chipselect),                             //                                               .chipselect
		.sram_s1_clken                                        (mm_interconnect_0_sram_s1_clken),                                  //                                               .clken
		.uart_avalon_jtag_slave_address                       (mm_interconnect_0_uart_avalon_jtag_slave_address),                 //                         uart_avalon_jtag_slave.address
		.uart_avalon_jtag_slave_write                         (mm_interconnect_0_uart_avalon_jtag_slave_write),                   //                                               .write
		.uart_avalon_jtag_slave_read                          (mm_interconnect_0_uart_avalon_jtag_slave_read),                    //                                               .read
		.uart_avalon_jtag_slave_readdata                      (mm_interconnect_0_uart_avalon_jtag_slave_readdata),                //                                               .readdata
		.uart_avalon_jtag_slave_writedata                     (mm_interconnect_0_uart_avalon_jtag_slave_writedata),               //                                               .writedata
		.uart_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest),             //                                               .waitrequest
		.uart_avalon_jtag_slave_chipselect                    (mm_interconnect_0_uart_avalon_jtag_slave_chipselect)               //                                               .chipselect
	);

	RedNeuronal_NiosII_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (redneuronal_niosii_irq_irq)      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (redneuronal_niosii_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),               // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),           //          .reset_req
		.reset_req_in0  (1'b0),                                         // (terminated)
		.reset_in1      (1'b0),                                         // (terminated)
		.reset_req_in1  (1'b0),                                         // (terminated)
		.reset_in2      (1'b0),                                         // (terminated)
		.reset_req_in2  (1'b0),                                         // (terminated)
		.reset_in3      (1'b0),                                         // (terminated)
		.reset_req_in3  (1'b0),                                         // (terminated)
		.reset_in4      (1'b0),                                         // (terminated)
		.reset_req_in4  (1'b0),                                         // (terminated)
		.reset_in5      (1'b0),                                         // (terminated)
		.reset_req_in5  (1'b0),                                         // (terminated)
		.reset_in6      (1'b0),                                         // (terminated)
		.reset_req_in6  (1'b0),                                         // (terminated)
		.reset_in7      (1'b0),                                         // (terminated)
		.reset_req_in7  (1'b0),                                         // (terminated)
		.reset_in8      (1'b0),                                         // (terminated)
		.reset_req_in8  (1'b0),                                         // (terminated)
		.reset_in9      (1'b0),                                         // (terminated)
		.reset_req_in9  (1'b0),                                         // (terminated)
		.reset_in10     (1'b0),                                         // (terminated)
		.reset_req_in10 (1'b0),                                         // (terminated)
		.reset_in11     (1'b0),                                         // (terminated)
		.reset_req_in11 (1'b0),                                         // (terminated)
		.reset_in12     (1'b0),                                         // (terminated)
		.reset_req_in12 (1'b0),                                         // (terminated)
		.reset_in13     (1'b0),                                         // (terminated)
		.reset_req_in13 (1'b0),                                         // (terminated)
		.reset_in14     (1'b0),                                         // (terminated)
		.reset_req_in14 (1'b0),                                         // (terminated)
		.reset_in15     (1'b0),                                         // (terminated)
		.reset_req_in15 (1'b0)                                          // (terminated)
	);

endmodule
