
module RedNeuronal_NiosII (
	clk_clk);	

	input		clk_clk;
endmodule
